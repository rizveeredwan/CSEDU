// DSCH3
// 4/24/2006 2:07:32 PM
// D:\Documents and Settings\AhsanReza\Desktop\NUB thesis\thesis presentations\vlsi simulator\dsch3\sajib.sym

module sajib( );
 wire w2,w3,w4,w5,w6;
 xor #(9) xor2_1(w4,w2,w3);
 xor #(16) xor2_2(w2,w5,w6);
endmodule

// Simulation parameters in Verilog Format

// Simulation parameters
